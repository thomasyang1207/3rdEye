library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Camera_Init is
	port(
		clk, rst: in std_logic;
		start: in std_logic;
		done: out std_logic;
		
		sda : inout std_logic; --serial data output of i2c bus
		scl : inout std_logic --serial clock output of i2c bus
	);
end Camera_Init;

architecture arch of Camera_Init is

	type state_type is (idle, sending, stop);
	
	signal state_reg: state_type := idle;
	signal state_next: state_type; 
	
	signal ind_reg: integer := 0;
	signal ind_next: integer;
	signal ind_succ: integer;
	
	type i2cframe is record
		addr: std_logic_vector(6 downto 0);
		rw: std_logic;
		write_one: std_logic; --1 if only register; 
		reg_wr: std_logic_vector(7 downto 0);
		data_wr: std_logic_vector(7 downto 0);
	end record;

	type i2cFrameArray is array(natural range<>) of i2cframe;
	
	constant initFile: i2cFrameArray := 
	(
		("0110000", '0', '0', x"ff", x"00"), 
		("0110000", '0', '0', x"2c", x"ff"), 
		("0110000", '0', '0', x"2e", x"df"), 
		("0110000", '0', '0', x"ff", x"01"), 
		("0110000", '0', '0', x"3c", x"32"), 
		("0110000", '0', '0', x"11", x"01"), 
		("0110000", '0', '0', x"09", x"02"), 
		("0110000", '0', '0', x"04", x"28"), 
		("0110000", '0', '0', x"13", x"e5"), 
		("0110000", '0', '0', x"14", x"48"), 
		("0110000", '0', '0', x"2c", x"0c"), 
		("0110000", '0', '0', x"33", x"78"), 
		("0110000", '0', '0', x"3a", x"33"), 
		("0110000", '0', '0', x"3b", x"fB"), 
		("0110000", '0', '0', x"3e", x"00"), 
		("0110000", '0', '0', x"43", x"11"), 
		("0110000", '0', '0', x"16", x"10"), 
		("0110000", '0', '0', x"39", x"92"), 
		("0110000", '0', '0', x"35", x"da"), 
		("0110000", '0', '0', x"22", x"1a"), 
		("0110000", '0', '0', x"37", x"c3"), 
		("0110000", '0', '0', x"23", x"00"), 
		("0110000", '0', '0', x"34", x"c0"), 
		("0110000", '0', '0', x"36", x"1a"), 
		("0110000", '0', '0', x"06", x"88"), 
		("0110000", '0', '0', x"07", x"c0"), 
		("0110000", '0', '0', x"0d", x"87"), 
		("0110000", '0', '0', x"0e", x"41"), 
		("0110000", '0', '0', x"4c", x"00"), 
		("0110000", '0', '0', x"48", x"00"), 
		("0110000", '0', '0', x"5B", x"00"), 
		("0110000", '0', '0', x"42", x"03"), 
		("0110000", '0', '0', x"4a", x"81"), 
		("0110000", '0', '0', x"21", x"99"), 
		("0110000", '0', '0', x"24", x"40"), 
		("0110000", '0', '0', x"25", x"38"), 
		("0110000", '0', '0', x"26", x"82"), 
		("0110000", '0', '0', x"5c", x"00"), 
		("0110000", '0', '0', x"63", x"00"), 
		("0110000", '0', '0', x"61", x"70"), 
		("0110000", '0', '0', x"62", x"80"), 
		("0110000", '0', '0', x"7c", x"05"), 
		("0110000", '0', '0', x"20", x"80"), 
		("0110000", '0', '0', x"28", x"30"), 
		("0110000", '0', '0', x"6c", x"00"), 
		("0110000", '0', '0', x"6d", x"80"), 
		("0110000", '0', '0', x"6e", x"00"), 
		("0110000", '0', '0', x"70", x"02"), 
		("0110000", '0', '0', x"71", x"94"), 
		("0110000", '0', '0', x"73", x"c1"), 
		("0110000", '0', '0', x"12", x"40"), 
		("0110000", '0', '0', x"17", x"11"), 
		("0110000", '0', '0', x"18", x"43"), 
		("0110000", '0', '0', x"19", x"00"), 
		("0110000", '0', '0', x"1a", x"4b"), 
		("0110000", '0', '0', x"32", x"09"), 
		("0110000", '0', '0', x"37", x"c0"), 
		("0110000", '0', '0', x"4f", x"60"), 
		("0110000", '0', '0', x"50", x"a8"), 
		("0110000", '0', '0', x"6d", x"00"), 
		("0110000", '0', '0', x"3d", x"38"), 
		("0110000", '0', '0', x"46", x"3f"), 
		("0110000", '0', '0', x"4f", x"60"), 
		("0110000", '0', '0', x"0c", x"3c"), 
		("0110000", '0', '0', x"ff", x"00"), 
		("0110000", '0', '0', x"e5", x"7f"), 
		("0110000", '0', '0', x"f9", x"c0"), 
		("0110000", '0', '0', x"41", x"24"), 
		("0110000", '0', '0', x"e0", x"14"), 
		("0110000", '0', '0', x"76", x"ff"), 
		("0110000", '0', '0', x"33", x"a0"), 
		("0110000", '0', '0', x"42", x"20"), 
		("0110000", '0', '0', x"43", x"18"), 
		("0110000", '0', '0', x"4c", x"00"), 
		("0110000", '0', '0', x"87", x"d5"), 
		("0110000", '0', '0', x"88", x"3f"), 
		("0110000", '0', '0', x"d7", x"03"), 
		("0110000", '0', '0', x"d9", x"10"), 
		("0110000", '0', '0', x"d3", x"82"), 
		("0110000", '0', '0', x"c8", x"08"), 
		("0110000", '0', '0', x"c9", x"80"), 
		("0110000", '0', '0', x"7c", x"00"), 
		("0110000", '0', '0', x"7d", x"00"), 
		("0110000", '0', '0', x"7c", x"03"), 
		("0110000", '0', '0', x"7d", x"48"), 
		("0110000", '0', '0', x"7d", x"48"), 
		("0110000", '0', '0', x"7c", x"08"), 
		("0110000", '0', '0', x"7d", x"20"), 
		("0110000", '0', '0', x"7d", x"10"), 
		("0110000", '0', '0', x"7d", x"0e"), 
		("0110000", '0', '0', x"90", x"00"), 
		("0110000", '0', '0', x"91", x"0e"), 
		("0110000", '0', '0', x"91", x"1a"), 
		("0110000", '0', '0', x"91", x"31"), 
		("0110000", '0', '0', x"91", x"5a"), 
		("0110000", '0', '0', x"91", x"69"), 
		("0110000", '0', '0', x"91", x"75"), 
		("0110000", '0', '0', x"91", x"7e"), 
		("0110000", '0', '0', x"91", x"88"), 
		("0110000", '0', '0', x"91", x"8f"), 
		("0110000", '0', '0', x"91", x"96"), 
		("0110000", '0', '0', x"91", x"a3"), 
		("0110000", '0', '0', x"91", x"af"), 
		("0110000", '0', '0', x"91", x"c4"), 
		("0110000", '0', '0', x"91", x"d7"), 
		("0110000", '0', '0', x"91", x"e8"), 
		("0110000", '0', '0', x"91", x"20"), 
		("0110000", '0', '0', x"92", x"00"), 
		("0110000", '0', '0', x"93", x"06"), 
		("0110000", '0', '0', x"93", x"e3"), 
		("0110000", '0', '0', x"93", x"05"), 
		("0110000", '0', '0', x"93", x"05"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"04"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"93", x"00"), 
		("0110000", '0', '0', x"96", x"00"), 
		("0110000", '0', '0', x"97", x"08"), 
		("0110000", '0', '0', x"97", x"19"), 
		("0110000", '0', '0', x"97", x"02"), 
		("0110000", '0', '0', x"97", x"0c"), 
		("0110000", '0', '0', x"97", x"24"), 
		("0110000", '0', '0', x"97", x"30"), 
		("0110000", '0', '0', x"97", x"28"), 
		("0110000", '0', '0', x"97", x"26"), 
		("0110000", '0', '0', x"97", x"02"), 
		("0110000", '0', '0', x"97", x"98"), 
		("0110000", '0', '0', x"97", x"80"), 
		("0110000", '0', '0', x"97", x"00"), 
		("0110000", '0', '0', x"97", x"00"), 
		("0110000", '0', '0', x"c3", x"ed"), 
		("0110000", '0', '0', x"a4", x"00"), 
		("0110000", '0', '0', x"a8", x"00"), 
		("0110000", '0', '0', x"c5", x"11"), 
		("0110000", '0', '0', x"c6", x"51"), 
		("0110000", '0', '0', x"bf", x"80"), 
		("0110000", '0', '0', x"c7", x"10"), 
		("0110000", '0', '0', x"b6", x"66"), 
		("0110000", '0', '0', x"b8", x"A5"), 
		("0110000", '0', '0', x"b7", x"64"), 
		("0110000", '0', '0', x"b9", x"7C"), 
		("0110000", '0', '0', x"b3", x"af"), 
		("0110000", '0', '0', x"b4", x"97"), 
		("0110000", '0', '0', x"b5", x"FF"), 
		("0110000", '0', '0', x"b0", x"C5"), 
		("0110000", '0', '0', x"b1", x"94"), 
		("0110000", '0', '0', x"b2", x"0f"), 
		("0110000", '0', '0', x"c4", x"5c"), 
		("0110000", '0', '0', x"c0", x"64"), 
		("0110000", '0', '0', x"c1", x"4B"), 
		("0110000", '0', '0', x"8c", x"00"), 
		("0110000", '0', '0', x"86", x"3D"), 
		("0110000", '0', '0', x"50", x"00"), 
		("0110000", '0', '0', x"51", x"C8"), 
		("0110000", '0', '0', x"52", x"96"), 
		("0110000", '0', '0', x"53", x"00"), 
		("0110000", '0', '0', x"54", x"00"), 
		("0110000", '0', '0', x"55", x"00"), 
		("0110000", '0', '0', x"5a", x"C8"), 
		("0110000", '0', '0', x"5b", x"96"), 
		("0110000", '0', '0', x"5c", x"00"), 
		("0110000", '0', '0', x"d3", x"00"), 
		("0110000", '0', '0', x"c3", x"ed"), 
		("0110000", '0', '0', x"7f", x"00"), 
		("0110000", '0', '0', x"da", x"00"), 
		("0110000", '0', '0', x"e5", x"1f"), 
		("0110000", '0', '0', x"e1", x"67"), 
		("0110000", '0', '0', x"e0", x"00"), 
		("0110000", '0', '0', x"dd", x"7f"), 
		("0110000", '0', '0', x"05", x"00"), 
		("0110000", '0', '0', x"12", x"40"), 
		("0110000", '0', '0', x"d3", x"04"), 
		("0110000", '0', '0', x"c0", x"16"), 
		("0110000", '0', '0', x"C1", x"12"), 
		("0110000", '0', '0', x"8c", x"00"), 
		("0110000", '0', '0', x"86", x"3d"), 
		("0110000", '0', '0', x"50", x"00"), 
		("0110000", '0', '0', x"51", x"2C"), 
		("0110000", '0', '0', x"52", x"24"), 
		("0110000", '0', '0', x"53", x"00"), 
		("0110000", '0', '0', x"54", x"00"), 
		("0110000", '0', '0', x"55", x"00"), 
		("0110000", '0', '0', x"5A", x"2c"), 
		("0110000", '0', '0', x"5b", x"24"), 
		("0110000", '0', '0', x"5c", x"00"), 
		("0110000", '0', '0', x"FF", x"00"), 
		("0110000", '0', '0', x"05", x"00"), 
		("0110000", '0', '0', x"DA", x"10"), 
		("0110000", '0', '0', x"D7", x"03"), 
		("0110000", '0', '0', x"DF", x"00"), 
		("0110000", '0', '0', x"33", x"80"), 
		("0110000", '0', '0', x"3C", x"40"), 
		("0110000", '0', '0', x"e1", x"77"), 
		("0110000", '0', '0', x"00", x"00"), 
		("0110000", '0', '0', x"e0", x"14"), 
		("0110000", '0', '0', x"e1", x"77"), 
		("0110000", '0', '0', x"e5", x"1f"), 
		("0110000", '0', '0', x"d7", x"03"), 
		("0110000", '0', '0', x"da", x"10"), 
		("0110000", '0', '0', x"e0", x"00"), 
		("0110000", '0', '0', x"FF", x"01"), 
		("0110000", '0', '0', x"04", x"08"), 
		("0110000", '0', '0', x"ff", x"01"), 
		("0110000", '0', '0', x"11", x"01"), 
		("0110000", '0', '0', x"12", x"00"), 
		("0110000", '0', '0', x"17", x"11"), 
		("0110000", '0', '0', x"18", x"75"), 
		("0110000", '0', '0', x"32", x"36"), 
		("0110000", '0', '0', x"19", x"01"), 
		("0110000", '0', '0', x"1a", x"97"), 
		("0110000", '0', '0', x"03", x"0f"), 
		("0110000", '0', '0', x"37", x"40"), 
		("0110000", '0', '0', x"4f", x"bb"), 
		("0110000", '0', '0', x"50", x"9c"), 
		("0110000", '0', '0', x"5a", x"57"), 
		("0110000", '0', '0', x"6d", x"80"), 
		("0110000", '0', '0', x"3d", x"34"), 
		("0110000", '0', '0', x"39", x"02"), 
		("0110000", '0', '0', x"35", x"88"), 
		("0110000", '0', '0', x"22", x"0a"), 
		("0110000", '0', '0', x"37", x"40"), 
		("0110000", '0', '0', x"34", x"a0"), 
		("0110000", '0', '0', x"06", x"02"), 
		("0110000", '0', '0', x"0d", x"b7"), 
		("0110000", '0', '0', x"0e", x"01"), 
		("0110000", '0', '0', x"ff", x"00"), 
		("0110000", '0', '0', x"e0", x"04"), 
		("0110000", '0', '0', x"c0", x"c8"), 
		("0110000", '0', '0', x"c1", x"96"), 
		("0110000", '0', '0', x"86", x"3d"), 
		("0110000", '0', '0', x"50", x"89"), 
		("0110000", '0', '0', x"51", x"90"), 
		("0110000", '0', '0', x"52", x"2c"), 
		("0110000", '0', '0', x"53", x"00"), 
		("0110000", '0', '0', x"54", x"00"), 
		("0110000", '0', '0', x"55", x"88"), 
		("0110000", '0', '0', x"57", x"00"), 
		("0110000", '0', '0', x"5a", x"a0"), 
		("0110000", '0', '0', x"5b", x"78"), 
		("0110000", '0', '0', x"5c", x"00"), 
		("0110000", '0', '0', x"d3", x"04"), 
		("0110000", '0', '0', x"e0", x"00")
	); 
	
	signal ena: std_logic;
	signal rw: std_logic;
	signal write_one: std_logic;
	signal slave_addr: std_logic_vector(6 downto 0);
	signal reg_wr: std_logic_vector(7 downto 0);
	signal data_wr: std_logic_vector(7 downto 0);
	signal data_rd: std_logic_vector(7 downto 0);
	signal done_transmit: std_logic;
	signal ready: std_logic;
	signal ack_error: std_logic;
	
	COMPONENT I2C
		port(
			clk : in std_logic; --system clock
			rst : in std_logic; --reset. Active HIGH reset. 
			ena : in std_logic; --enable => assert 1 when the data is ready. Don't assert if you don't want the system to leave idle mode.
			
			rw : in std_logic; --0 is write; 1 is read. good to use something like addr & rw
			write_one: in std_logic; --1 to write only the register, 0 to write both register and data. 
			
			slave_addr: in std_logic_vector(6 downto 0); --7-bit address, for our application, it will be 0x30
			reg_wr: in std_logic_vector(7 downto 0); 
			data_wr : in std_logic_vector(7 downto 0); --data to write to slave;
		
			data_rd : out STD_LOGIC_VECTOR(7 downto 0); --data read from slave
			
			done_transmit : out std_logic; --single pulse indicating that the data_rd is valid
			ready: out std_logic; --signal indicating that the device is ready. 
			ack_error : out std_logic; --flag if improper acknowledge from slave; i.e. if slave was reset, etc.
			
			sda : inout std_logic; --serial data output of i2c bus
			scl : inout std_logic --serial clock output of i2c bus
		);
	end COMPONENT;

begin
	I2c_inst: I2C port map(clk => clk, rst => rst, ena => ena, rw => rw,
								  write_one => write_one, slave_addr => slave_addr, reg_wr => reg_wr,
								  data_wr => data_wr, data_rd => data_rd, done_transmit => done_transmit,
								  ready => ready, ack_error => ack_error, sda => sda, scl => scl);
	
	
	
	slave_addr <= initFile(ind_reg).addr;
	rw <= initFile(ind_reg).rw;
	write_one <= initFile(ind_reg).write_one;
	reg_wr <= initFile(ind_reg).reg_Wr;
	data_wr <= initFile(ind_reg).data_wr;
	
	ind_succ <= ind_reg + 1;
	
	clocked: process(clk, rst)
	begin
		if rst = '1' then
			state_reg <= idle;
			ind_reg <= 0;
		elsif rising_edge(clk) then
			state_reg <= state_next;
			ind_reg <= ind_next;
		end if;
	end process;
	
	get_next: process(state_reg, ind_reg, start, ready, ind_succ, done_transmit, ack_error)
	begin
		state_next <= state_reg;
		ind_next <= ind_reg;
		ena <= '0';
		done <= '0';
		
		case state_reg is
			when idle =>
				if start = '1' then
					state_next <= sending;
					ind_next <= 0;
				end if;
			when sending => 
				--if the i2c isn't sending anything right now, send an enable signal, and then update the i2c...
				if ready = '1' then
					ena <= '1'; --begin to start...
				end if;
				
				if done_transmit = '1' then
					--time to increment stuff...
					if ind_succ < initFile'length then
						ind_next <= ind_succ;
					else
						state_next <= stop;
					end if;
				end if;
				
				if ack_error = '1' then
					ind_next <= 0;
				end if;
			
			when stop => 
				done <= '1';
				state_next <= idle;
				
			when others =>
		end case;
	
	end process;

end arch;