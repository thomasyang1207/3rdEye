--Webcam; topmost entity; 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Webcam is
	port(
		-- Camera ports
		Data_bus: in std_logic_vector(7 downto 0);	
		pclk: in std_logic;
		href: in std_logic; 
		vsync: in std_logic; 
		
		
		xclk: out std_logic; 
		sda: inout std_logic; 
		scl: out std_logic; 
		rst: out std_logic; 
		
		
		--SRAM Ports 
		sram_addr: out std_logic_vector(19 downto 0); 
		sram_data: inout std_logic_vector(15 downto 0);
		we_sram: out std_logic; -- output 
		oe_sram: out std_logic; --output enable; assert 0 to read
		
		ce: out std_logic; 
		ub: out std_logic; 
		lb: out std_logic; 
		
		
		
		--display ports
		digit1, digit2, digit3, digit4: out std_logic_vector(6 downto 0); 
		
		
		
		--read pins 
		read_on: in std_logic; 
		
		--general
		clk: in std_logic 
	
	);
end Webcam;



architecture arch of Webcam is

	COMPONENT camera_controller
		PORT(
			-- interface with the main system; 
			clk    : in    STD_LOGIC;
			resend : in    STD_LOGIC; -- by default, we begin the resend pin set high; 
			config_finished : out std_logic;
	 
		-- interface with camera; 
			sioc  : out   STD_LOGIC; -- provided TO the OV2640; 
			siod  : inout STD_LOGIC; -- i2c data wire; 
		
			-- hold these constant; 
			reset : out   STD_LOGIC; -- reset signal to the camera;
			xclk  : out   STD_LOGIC
		);
	end COMPONENT; 
	
	
	
	COMPONENT parallel_capture
		PORT(
			--from camera: 
			pclk: in std_logic;
			href: in std_logic;
			vsync: in std_logic; 
			data_bus: in std_logic_vector(7 downto 0); 
			
			--from fpga (central unit): 
			read_i: in std_logic; -- signal to BE in read process; -- do we need this? 
			
			--to FPGA (SRAM controller)
			we_o: out std_logic; -- always 0; 
			mem_o: out std_logic; 
			addr_o: out std_logic_vector(19 downto 0); --generated by the address generator; 
			data_o: out std_logic_vector(15 downto 0); --think about the design here; 
			
			image_available_out: out std_logic
		);
	end COMPONENT;
	
	COMPONENT sram_controller
		PORT(
			addr_i: in std_logic_vector(19 downto 0); --20 bit address; 
			data_i: in std_logic_vector(15 downto 0); 
			we_i: in std_logic; 
			mem_i: in std_logic; 
			
			--outputs from interface
			data_o: out std_logic_vector(15 downto 0);
			ready: out std_logic; 
			
			--inputs to sram
			sram_addr_o: out std_logic_vector(19 downto 0); 
			sram_data_io: inout std_logic_vector(15 downto 0);
			we_o: out std_logic; -- output 
			oe_o: out std_logic; --output enable; assert 0 to read
		
		
			--clk and reset: 
			clk_i, reset_i: in std_logic
		);
	end COMPONENT;
	
	
	COMPONENT control_unit 
		PORT(
			--general signals:
			clk: in std_logic; 
		
			--from i2c sender; 
			resend_init: out std_logic; 
			camera_config_finished: in std_logic; 
		
			--camera reader: 
			image_available: in std_logic; -- just a signal that is set high when image has finished transferring. 
			capture_on: out std_logic; 
			
			--address selection
			select_signal: out std_logic;
		
			--demo portion 
			read_on: in std_logic -- how to enter read mode; 
			--UART control - coming soon! 
		);
	end COMPONENT;
	
	COMPONENT rw_mux
		PORT(
			select_i: in std_logic; -- selects the data; 
			addr1_i: in std_logic_vector(19 downto 0);
			we1_i: in std_logic; 
			mem1_i: in std_logic; 
			
			addr2_i: in std_logic_vector(19 downto 0);
			we2_i: in std_logic; 
			mem2_i: in std_logic; 
			
			we_o: out std_logic; 
			mem_o: out std_logic; 
			addr_o: out std_logic_vector(19 downto 0)
		);
	end COMPONENT;
	
	
	
	COMPONENT LED_converter 
		PORT(
			in1: in std_logic_vector(3 downto 0); 
			out1: out std_logic_vector(6 downto 0)
		);
	end COMPONENT; 
	
	

	signal display_reg: std_logic_vector(15 downto 0) := x"43a2"; 
	signal read_addr: std_logic_vector(19 downto 0) := (others => '0'); 
	
	--internal signals! 
	signal camera_resend: std_logic; 
	signal camera_config_finished: std_logic; 
	
	signal image_available: std_logic; 
	signal capture_on: std_logic;
	
	signal rw_mux_select: std_logic; 
	
	
	signal addr1: std_logic_vector(19 downto 0);
	signal addr2: std_logic_vector(19 downto 0);	
	signal addr_out: std_logic_vector(19 downto 0);
	
	signal we1: std_logic;
	signal we2: std_logic;	
	signal we_out: std_logic;
	
	signal mem1: std_logic;
	signal mem2: std_logic;	
	signal mem_out: std_logic;
	
	signal data_in: std_logic_vector(15 downto 0); -- data into the SRAM, 
	signal data_out: std_logic_vector(15 downto 0); -- data coming out of the sram; 
	signal sram_reset: std_logic := '0'; 
	
	
	
	--SRAM READS 
	signal sram_ready: std_logic;

begin
	
	camera_controller_inst: camera_controller port map(
		clk => clk, 
		resend => camera_resend,
		config_finished => camera_config_finished,
		sioc => scl, 
		siod => sda, 
		reset => rst, 
		xclk => xclk
	); 
	
	
	
	parallel_capture_inst: parallel_capture port map(
		pclk => pclk, 
		href => href, 
		vsync => vsync, 
		data_bus => Data_bus,
		
		read_i => capture_on, 
		
		we_o => we1, 
		mem_o => mem1, 
		addr_o => addr1, 
		data_o => data_in,
		
		image_available_out => image_available
	);

	
	
	
	sram_controller_inst: sram_controller port map(
		addr_i => addr_out, 
		data_i => data_in, 
		we_i => we_out,
		mem_i => mem_out, 
		
		--outputs from interface
		data_o => data_out, 
		ready => sram_ready,
		
		--inputs to sram
		sram_addr_o => sram_addr, 
		sram_data_io => sram_data,
		we_o => we_sram, -- output 
		oe_o => oe_sram, --output enable; assert 0 to read
		
		
		--clk and reset: 
		clk_i => clk,
		reset_i => sram_reset
	);
	
	
	
	
	control_unit_inst: control_unit port map(
		clk => clk, 
		resend_init => camera_resend, 
		camera_config_finished => camera_config_finished, 
		
		image_available => image_available, 
		capture_on => capture_on, 
		select_signal => rw_mux_select, 
		
		read_on => read_on 
	); 
	
	
	rw_mux_inst: rw_mux port map(
		select_i => rw_mux_select, 
		addr1_i => addr1, 
		we1_i => we1, 
		mem1_i => mem1,  
		
		addr2_i => addr2, 
		we2_i => we2, 
		mem2_i => mem2, 
		
		we_o => we_out, 
		mem_o => mem_out,
		addr_o => addr_out 
	); 
	
	LED1: LED_converter port map(
		in1 => display_reg(11 downto 8), 
		out1 => digit1
	);
	
	LED2: LED_converter port map(
		in1 => display_reg(15 downto 12),
		out1 => digit2
	);
	
	LED3: LED_converter port map(
		in1 => display_reg(3 downto 0), 
		out1 => digit3
	);
	
	LED4: LED_converter port map(
		in1 => display_reg(7 downto 4), 
		out1 => digit4
	);
	
	process(clk, mem_out, rw_mux_select) -- process to set the display register, when we have an output read. 
	begin 
		if rising_edge(clk) then
					display_reg <= data_out; -- read mode register;
		end if; 
	end process; 

	
	ce <= '0';  
	ub <= '0';  
	lb <= '0'; 
	

end arch; 