library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity parallel_capture is
	port(
		--from camera: 
		pclk: in std_logic;
		href: in std_logic;
		vsync: in std_logic; 
		data_bus: in std_logic_vector(7 downto 0); 
		
		--from fpga (central unit): 
		read_i: in std_logic; -- signal to BE in read process; -- do we need this? 
		
		--to FPGA (SRAM controller)
		we_o: out std_logic; -- always 0; 
		mem_o: out std_logic; 
		addr_o: out std_logic_vector(19 downto 0); --generated by the address generator; 
		data_o: out std_logic_vector(15 downto 0); --think about the design here; 
		
		image_available_out: out std_logic
		
	); 
end parallel_capture; 


architecture arch of parallel_capture is 
	
	Component address_generator 
	port(
	
		new_addr: in std_logic; -- set to 1, to enable new address to be written; basically the reset signal; 
		advance_addr: in std_logic; -- only increment the address when this is set high 
		
		clk: in std_logic; -- pclk; 
		addr: out std_logic_vector(19 downto 0) --19 bit address here; 
	);
	end component;
	
	
	--signals and registers; 
	signal ffd8: std_logic; 
	signal advance: std_logic; -- don't advance if we didn't actually receive 
	signal advance_next: std_logic; -- don't advance if we didn't actually receive 
	signal mem_r: std_logic; 
	signal mem_next: std_logic; 
	
	--data registers 
	signal data_reg1: std_logic_vector(7 downto 0); 
	signal data_reg2: std_logic_vector(7 downto 0); -- map these into the outputs; --write every 
	
	--hsync and vref states; 
	type capture_state_type is (wait1, wait2, capture1, capture2, done1, done2); --capture 1-> capture and write on, capture 2-> capture and write OFF; 
	signal capture_state: capture_state_type;
	signal capture_state_next: capture_state_type; 
	
	signal image_available: std_logic; 
	
	
begin
	--default values 
	we_o <= '0'; -- write; 
	ffd8 <= '1' when (data_reg1 = x"FF" and data_bus = x"D8") else '0'; 
	image_available <= '1' when (data_reg2 = x"FF" and data_reg1 = x"D9") else '0'; --
	
	--clocked
	process(pclk, vsync, read_i)
	begin
		if rising_edge(pclk) then
				data_reg2 <= data_reg1; 
				if(vsync = '1') then
					data_reg1 <= data_bus;
				else 
					data_reg1 <= (others => '0'); -- if there isn't a new byte, then we will go to 0. 
				end if; 
				capture_state <= capture_state_next; 
				advance <= advance_next; 
				mem_r <= mem_next; 
		end if;
	end process; 
	
	--unclocked
	
	process(capture_state_next, vsync, href)
	begin 
		image_available_out <= '0'; 
		case capture_state_next is 
			when wait1 => 
				advance_next <= '0'; 
				mem_next <= '0'; 
			
			when wait2 =>
				advance_next <= '0'; 
				mem_next <= '0'; 
			
			when capture1 =>
				advance_next <= '0'; 
				mem_next <= '0'; 
			
			when capture2 =>
				advance_next <= '1'; -- retrieve NEW address on NEXT clock cycle;  
				mem_next <= '1'; --capture only HERE; 
				
			when done1 => 
				advance_next <= '0'; 
				mem_next <= '0'; -- stay here until we receive another read request; 
				image_available_out <= '1'; 
				
			when done2 => 
				advance_next <= '0'; 
				mem_next <= '0'; 
				image_available_out <= '1'; 
		end case; 
	
	end process;
	
		--next state: 
	process(capture_state, vsync, href, ffd8, image_available, read_i)
	begin 
		--default 
		
		--other 
		case capture_state is 
			when wait1 => 
				capture_state_next <= wait1; --default; 
				--unless vsync is HIGH
				if(vsync = '1') then
					capture_state_next <= wait2; 
				end if; 
			
			
			when wait2 => 
				capture_state_next <= wait2; 
				if (vsync = '0') then 
					capture_state_next <= wait1; 
				elsif (ffd8 = '1') then
					capture_state_next <= capture1; 
				end if; 
			
			when capture1 => 
				capture_state_next <= capture2; --must go to the second capture state, regardless of whether capture has ended; 
			
			when capture2 => 
				capture_state_next <= capture2; 
				if (vsync = '0' and href = '0') then
					capture_state_next <= done1; 
				elsif (image_available = '1') then
					capture_state_next <= done1; 
				elsif (vsync = '0') then 
					capture_state_next <= done1; 
				end if; 
			
			when done1 => 
				capture_state_next <= done2; 
				
				
			when done2 => 
				capture_state_next <= done2; 
				if(read_i = '1') then 
					capture_state_next <= wait1; --effectively resetting the state; 
				end if; 
		
		end case; 
	
	end process; 
	
	
	--component maps: 
	addr_gen_inst: address_generator port map(
		new_addr => ffd8, -- new addr - set if the incoming byte is ffd8; 
		advance_addr => advance, --advance 
		clk => pclk, 
		addr => addr_o
	); 
	
	
	--outputs: 
	mem_o <= mem_r; 
	data_o <= data_reg1 & data_reg2; 

end arch; 